`ifndef EXECUTE_TYPES_SVH
`define EXECUTE_TYPES_SVH

package execute_types;
    typedef struct packed {logic clk;} input_t;

    typedef struct packed {logic clk;} output_t;
endpackage

`endif
